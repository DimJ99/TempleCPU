// #include 
/////////////////////////////////////////////////////////////////////////////////////////
/*
Contributor(s):


Parameter Descriptions:


*/
/////////////////////////////////////////////////////////////////////////////////////////


module insert_name 

// #(

// )

(
    input logic clk, n_rst
);


endmodule

/////////////////////////////////////////////////////////////////////////////////////////
/*
Sources (If deemed necessary, otherwise remove section):
(Just a link)

*/
/////////////////////////////////////////////////////////////////////////////////////////
